package pkg;


	
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "ahb_xtn.sv"
	`include "ahb_config.sv"
	`include "apb_config.sv"
	`include "env_config.sv"
	`include "ahb_drv.sv"
	`include "ahb_mon.sv"
	`include "ahb_seqr.sv"
	`include "ahb_agt.sv"
	`include "ahb_top.sv"
	`include "ahb_seq.sv"

	`include "apb_xtn.sv"
	`include "apb_mon.sv"
	`include "apb_seqr.sv"
	`include "apb_seq.sv"

	`include "apb_drv.sv"

	//`include "apb_seq.sv"
	`include "apb_agt.sv"
	`include "apb_top.sv"

	`include "virtual_seqr.sv"
	`include "virtual_seqs.sv"
	`include "scoreboard.sv"

	`include "tb.sv"


	`include "vtest.sv"
	
endpackage
